`default_nettype none

module top(input i_clock);
    always @ (posedge i_clock)
    begin
    end
endmodule
